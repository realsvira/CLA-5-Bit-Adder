magic
tech scmos
timestamp 1731580654
<< nwell >>
rect 28 -189 114 -90
rect 28 -208 126 -189
rect 100 -229 126 -208
<< ntransistor >>
rect 112 -252 114 -242
rect 39 -264 41 -254
rect 51 -264 53 -254
rect 63 -264 65 -254
rect 75 -264 77 -254
rect 87 -264 89 -254
<< ptransistor >>
rect 39 -202 41 -102
rect 51 -202 53 -102
rect 63 -202 65 -102
rect 75 -202 77 -102
rect 87 -202 89 -102
rect 112 -222 114 -202
<< ndiffusion >>
rect 111 -252 112 -242
rect 114 -252 115 -242
rect 38 -264 39 -254
rect 41 -264 42 -254
rect 50 -264 51 -254
rect 53 -264 54 -254
rect 62 -264 63 -254
rect 65 -264 66 -254
rect 74 -264 75 -254
rect 77 -264 78 -254
rect 86 -264 87 -254
rect 89 -264 90 -254
<< pdiffusion >>
rect 38 -202 39 -102
rect 41 -202 51 -102
rect 53 -202 63 -102
rect 65 -202 75 -102
rect 77 -202 87 -102
rect 89 -202 90 -102
rect 111 -222 112 -202
rect 114 -222 115 -202
<< ndcontact >>
rect 107 -252 111 -242
rect 115 -252 119 -242
rect 34 -264 38 -254
rect 42 -264 50 -254
rect 54 -264 62 -254
rect 66 -264 74 -254
rect 78 -264 86 -254
rect 90 -264 94 -254
<< pdcontact >>
rect 34 -202 38 -102
rect 90 -202 94 -102
rect 107 -222 111 -202
rect 115 -222 119 -202
<< psubstratepcontact >>
rect 107 -264 111 -260
rect 34 -273 38 -269
rect 44 -273 48 -269
rect 56 -273 60 -269
rect 68 -273 72 -269
rect 80 -273 84 -269
rect 90 -273 94 -269
<< nsubstratencontact >>
rect 34 -97 38 -93
rect 43 -97 47 -93
rect 55 -97 59 -93
rect 67 -97 71 -93
rect 79 -97 83 -93
rect 89 -97 93 -93
rect 107 -194 111 -189
<< polysilicon >>
rect 39 -102 41 -99
rect 51 -102 53 -99
rect 63 -102 65 -99
rect 75 -102 77 -99
rect 87 -102 89 -99
rect 112 -202 114 -199
rect 39 -254 41 -202
rect 51 -254 53 -202
rect 63 -254 65 -202
rect 75 -254 77 -202
rect 87 -254 89 -202
rect 112 -242 114 -222
rect 112 -257 114 -252
rect 39 -267 41 -264
rect 51 -267 53 -264
rect 63 -267 65 -264
rect 75 -267 77 -264
rect 87 -267 89 -264
<< polycontact >>
rect 35 -215 39 -211
rect 47 -222 51 -218
rect 59 -229 63 -225
rect 71 -236 75 -232
rect 83 -243 87 -239
rect 108 -237 112 -233
<< metal1 >>
rect 34 -93 111 -92
rect 38 -97 43 -93
rect 47 -97 55 -93
rect 59 -97 67 -93
rect 71 -97 79 -93
rect 83 -97 89 -93
rect 93 -97 111 -93
rect 34 -98 111 -97
rect 34 -102 38 -98
rect 28 -215 35 -211
rect 28 -222 47 -218
rect 28 -229 59 -225
rect 28 -236 71 -232
rect 90 -233 94 -202
rect 107 -189 111 -98
rect 107 -202 111 -194
rect 115 -233 119 -222
rect 90 -237 108 -233
rect 115 -237 126 -233
rect 28 -243 83 -239
rect 90 -246 94 -237
rect 115 -242 119 -237
rect 42 -251 94 -246
rect 42 -254 50 -251
rect 66 -254 74 -251
rect 90 -254 94 -251
rect 107 -260 111 -252
rect 34 -268 38 -264
rect 54 -268 62 -264
rect 78 -268 86 -264
rect 107 -268 111 -264
rect 34 -269 111 -268
rect 38 -273 44 -269
rect 48 -273 56 -269
rect 60 -273 68 -269
rect 72 -273 80 -269
rect 84 -273 90 -269
rect 94 -273 111 -269
<< labels >>
rlabel metal1 62 -272 65 -270 1 gnd
rlabel metal1 30 -242 33 -240 3 a
rlabel metal1 30 -235 33 -233 3 b
rlabel metal1 30 -228 33 -226 3 c
rlabel metal1 30 -221 33 -219 3 d
rlabel metal1 30 -214 33 -212 3 e
rlabel metal1 62 -96 65 -94 5 vdd
rlabel metal1 121 -235 126 -234 7 out
rlabel metal1 91 -236 93 -234 1 nout
<< end >>
