* Saumya 2024102044

.include TSMC_180nm.txt
.param SUPPLY=1.8
.option scale=90n
.global gnd vdd

Vdd vdd gnd 'SUPPLY'

.option scale=0.09u

M1000 nout d vdd vdd CMOSP w=20 l=2
+  ad=400 pd=120 as=500 ps=210
M1001 vdd a nout vdd CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 out nout vdd vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1003 vdd c nout vdd CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 a_0_n84# c a_n12_n84# Gnd CMOSN w=40 l=2
+  ad=400 pd=100 as=400 ps=100
M1005 a_12_n84# b a_0_n84# Gnd CMOSN w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1006 nout a a_12_n84# Gnd CMOSN w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1007 a_n12_n84# d gnd Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=250 ps=120
M1008 out nout gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1009 nout b vdd vdd CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
C0 b c 0.42fF
C1 c a 0.08fF
C2 b a 0.59fF
C3 d nout 0.05fF
C4 c nout 0.20fF
C5 b nout 0.08fF
C6 nout out 0.05fF
C7 nout a 0.13fF
C8 d vdd 0.07fF
C9 gnd out 0.13fF
C10 c vdd 0.07fF
C11 gnd a 0.05fF
C12 b vdd 0.07fF
C13 out vdd 0.29fF
C14 vdd a 0.07fF
C15 gnd nout 0.47fF
C16 d c 0.26fF
C17 b d 0.08fF
C18 nout vdd 1.09fF
C19 d a 0.08fF
C20 gnd Gnd 0.49fF
C21 out Gnd 0.07fF
C22 nout Gnd 0.40fF
C23 a Gnd 0.37fF
C24 b Gnd 0.34fF
C25 c Gnd 0.30fF
C26 d Gnd 0.27fF
C27 vdd Gnd 3.57fF

va a gnd pulse 0 1.8 0 0.1n 0.1n 5n 10n
vb b gnd pulse 0 1.8 0 0.1n 0.1n 10n 20n
vc c gnd pulse 0 1.8 0 0.1n 0.1n 20n 40n
vd d gnd pulse 0 1.8 0 0.1n 0.1n 40n 80n
.tran 0.01n 120n

.control
run
set hcopypscolor = 1
set color0 = white   
set color1 = black   
plot v(a) v(b)+2 v(c)+4 v(d)+6 v(out)+8
set hcopypscolor = 1
set color0=white
set color1=black
.endc