* Saumya 2024102044
.include TSMC_180nm.txt
.param SUPPLY=1.8
.option scale=90n
.global gnd vdd

Vdd vdd gnd 'SUPPLY'
.option scale=0.09u

M1000 nout b vdd w_n22_n17# CMOSP w=20 l=2
+  ad=200 pd=60 as=364 ps=214
M1001 out nout gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=214 ps=144
M1002 out nout vdd w_n22_n17# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1003 vdd a nout w_n22_n17# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 a_n9_n56# b gnd Gnd CMOSN w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1005 nout a a_n9_n56# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
C0 out gnd 0.13fF
C1 a nout 0.19fF
C2 vdd out 0.23fF
C3 nout w_n22_n17# 0.11fF
C4 nout b 0.04fF
C5 a w_n22_n17# 0.07fF
C6 a b 0.19fF
C7 w_n22_n17# b 0.07fF
C8 nout gnd 0.07fF
C9 a gnd 0.04fF
C10 nout out 0.05fF
C11 vdd nout 0.50fF
C12 out w_n22_n17# 0.05fF
C13 vdd w_n22_n17# 0.34fF
C14 gnd Gnd 0.33fF
C15 out Gnd 0.08fF
C16 nout Gnd 0.31fF
C17 a Gnd 0.26fF
C18 b Gnd 0.22fF
C19 vdd Gnd 0.01fF
C20 w_n22_n17# Gnd 2.43fF

va a gnd pulse 0 1.8 0 0.1n 0.1n 10n 20n
vb b gnd pulse 0 1.8 0 0.1n 0.1n 20n 40n

.tran  0.01n 100ns
.control
run
set hcopypscolor = 1
set color0 = white   
set color1 = black   
plot v(a) v(b)+2 v(out)+4 title 'Saumya 2024102044'
set hcopypscolor = 1
set color0=white
set color1=black
.endc