magic
tech scmos
timestamp 1731575492
<< nwell >>
rect -40 -18 46 79
<< ntransistor >>
rect 32 -41 34 -31
rect -29 -61 -27 -51
rect -17 -61 -15 -51
rect -5 -61 -3 -51
rect 7 -61 9 -51
<< ptransistor >>
rect -29 -12 -27 68
rect -17 -12 -15 68
rect -5 -12 -3 68
rect 7 -12 9 68
rect 32 -11 34 9
<< ndiffusion >>
rect 31 -41 32 -31
rect 34 -41 35 -31
rect -30 -61 -29 -51
rect -27 -61 -26 -51
rect -18 -61 -17 -51
rect -15 -61 -14 -51
rect -6 -61 -5 -51
rect -3 -61 -2 -51
rect 6 -61 7 -51
rect 9 -61 10 -51
<< pdiffusion >>
rect -30 -12 -29 68
rect -27 -12 -17 68
rect -15 -12 -5 68
rect -3 -12 7 68
rect 9 -12 10 68
rect 31 -11 32 9
rect 34 -11 35 9
<< ndcontact >>
rect 27 -41 31 -31
rect 35 -41 39 -31
rect -34 -61 -30 -51
rect -26 -61 -18 -51
rect -14 -61 -6 -51
rect -2 -61 6 -51
rect 10 -61 14 -51
<< pdcontact >>
rect -34 -12 -30 68
rect 10 -12 14 68
rect 27 -11 31 9
rect 35 -11 39 9
<< psubstratepcontact >>
rect 27 -55 31 -51
rect -34 -69 -30 -65
rect -24 -69 -20 -65
rect -12 -69 -8 -65
rect 0 -69 4 -65
rect 10 -69 14 -65
<< nsubstratencontact >>
rect -34 72 -30 76
rect -25 72 -21 76
rect -13 72 -9 76
rect 0 72 4 76
rect 10 72 14 76
rect 27 15 31 19
<< polysilicon >>
rect -29 68 -27 71
rect -17 68 -15 71
rect -5 68 -3 71
rect 7 68 9 71
rect 32 9 34 12
rect -29 -51 -27 -12
rect -17 -51 -15 -12
rect -5 -51 -3 -12
rect 7 -51 9 -12
rect 32 -31 34 -11
rect 32 -46 34 -41
rect -29 -64 -27 -61
rect -17 -64 -15 -61
rect -5 -64 -3 -61
rect 7 -64 9 -61
<< polycontact >>
rect -34 -46 -29 -42
rect -22 -39 -17 -35
rect -10 -32 -5 -28
rect 2 -25 7 -21
rect 28 -26 32 -22
<< metal1 >>
rect -30 72 -25 76
rect -21 72 -13 76
rect -9 72 0 76
rect 4 72 10 76
rect 14 72 31 76
rect -34 68 -30 72
rect 27 19 31 72
rect 31 15 45 19
rect 27 9 31 15
rect -40 -25 2 -21
rect 10 -22 14 -12
rect 35 -22 39 -11
rect 10 -26 28 -22
rect 35 -26 46 -22
rect -40 -32 -10 -28
rect -40 -39 -22 -35
rect 10 -42 14 -26
rect 35 -31 39 -26
rect -40 -46 -34 -42
rect -26 -48 14 -42
rect -26 -51 -18 -48
rect -2 -51 6 -48
rect 27 -51 31 -41
rect -34 -65 -30 -61
rect -14 -65 -6 -61
rect 10 -65 14 -61
rect 27 -65 31 -55
rect -30 -69 -24 -65
rect -20 -69 -12 -65
rect -8 -69 0 -65
rect 4 -69 10 -65
rect 14 -69 31 -65
<< labels >>
rlabel metal1 -39 -45 -37 -43 3 a
rlabel metal1 -39 -38 -37 -36 3 b
rlabel metal1 -39 -31 -37 -29 3 c
rlabel metal1 -39 -24 -37 -22 3 d
rlabel metal1 -7 73 -5 75 5 vdd
rlabel metal1 -6 -68 -4 -66 1 gnd
rlabel metal1 41 -24 46 -23 7 out
rlabel metal1 12 -25 14 -23 1 nout
<< end >>
