magic
tech scmos
timestamp 1731574387
<< nwell >>
rect -22 -26 52 48
rect -22 -29 26 -26
<< ntransistor >>
rect 38 -49 40 -39
rect -11 -69 -9 -59
rect 1 -69 3 -59
rect 13 -69 15 -59
<< ptransistor >>
rect -11 -23 -9 37
rect 1 -23 3 37
rect 13 -23 15 37
rect 38 -19 40 1
<< ndiffusion >>
rect 37 -49 38 -39
rect 40 -49 41 -39
rect -12 -69 -11 -59
rect -9 -69 -8 -59
rect 0 -69 1 -59
rect 3 -69 4 -59
rect 12 -69 13 -59
rect 15 -69 16 -59
<< pdiffusion >>
rect -12 -23 -11 37
rect -9 -23 1 37
rect 3 -23 13 37
rect 15 -23 16 37
rect 37 -19 38 1
rect 40 -19 41 1
<< ndcontact >>
rect 33 -49 37 -39
rect 41 -49 45 -39
rect -16 -69 -12 -59
rect -8 -69 0 -59
rect 4 -69 12 -59
rect 16 -69 20 -59
<< pdcontact >>
rect -16 -23 -12 37
rect 16 -23 20 37
rect 33 -19 37 1
rect 41 -19 45 1
<< psubstratepcontact >>
rect -16 -79 -12 -75
rect -6 -79 -2 -75
rect 6 -79 10 -75
rect 16 -79 20 -75
<< nsubstratencontact >>
rect -16 41 -12 45
rect -7 41 -3 45
rect 5 41 9 45
rect 16 41 20 45
<< polysilicon >>
rect -11 37 -9 40
rect 1 37 3 40
rect 13 37 15 40
rect 38 1 40 4
rect -11 -59 -9 -23
rect 1 -59 3 -23
rect 13 -59 15 -23
rect 38 -39 40 -19
rect 38 -54 40 -49
rect -11 -72 -9 -69
rect 1 -72 3 -69
rect 13 -72 15 -69
<< polycontact >>
rect -16 -35 -11 -31
rect -4 -42 1 -38
rect 8 -49 13 -45
rect 34 -34 38 -30
<< metal1 >>
rect -12 41 -7 45
rect -3 41 5 45
rect 9 41 16 45
rect 20 41 37 45
rect -16 37 -12 41
rect 33 1 37 41
rect 16 -30 20 -23
rect 41 -30 45 -19
rect -22 -35 -16 -31
rect 16 -34 34 -30
rect 41 -34 52 -30
rect -22 -42 -4 -38
rect -22 -49 8 -45
rect 16 -52 20 -34
rect 41 -39 45 -34
rect -8 -56 20 -52
rect -8 -59 0 -56
rect 16 -59 20 -56
rect 33 -55 37 -49
rect 33 -59 45 -55
rect -16 -74 -12 -69
rect 4 -74 12 -69
rect -16 -75 20 -74
rect -12 -79 -6 -75
rect -2 -79 6 -75
rect 10 -79 16 -75
<< labels >>
rlabel metal1 -22 -48 -20 -46 3 c
rlabel metal1 -21 -41 -19 -39 3 b
rlabel metal1 -21 -34 -19 -32 3 a
rlabel metal1 47 -32 52 -31 7 out
rlabel metal1 36 -58 41 -57 1 gnd
rlabel metal1 -1 42 2 44 5 vdd
rlabel metal1 17 -33 19 -31 1 nout
rlabel metal1 0 -78 2 -76 1 gnd
<< end >>
