magic
tech scmos
timestamp 1764443331
<< nwell >>
rect -23 -17 49 26
<< ntransistor >>
rect 35 -37 37 -27
rect -12 -71 -10 -41
rect 0 -71 2 -41
rect 12 -71 14 -41
<< ptransistor >>
rect -12 -11 -10 9
rect 0 -11 2 9
rect 12 -11 14 9
rect 35 -7 37 13
<< ndiffusion >>
rect 34 -37 35 -27
rect 37 -37 38 -27
rect -13 -71 -12 -41
rect -10 -71 0 -41
rect 2 -71 12 -41
rect 14 -71 15 -41
<< pdiffusion >>
rect -13 -11 -12 9
rect -10 -11 -9 9
rect -1 -11 0 9
rect 2 -11 3 9
rect 11 -11 12 9
rect 14 -11 15 9
rect 34 -7 35 13
rect 37 -7 38 13
<< ndcontact >>
rect 30 -37 34 -27
rect 38 -37 42 -27
rect -17 -71 -13 -41
rect 15 -71 19 -41
<< pdcontact >>
rect -17 -11 -13 9
rect -9 -11 -1 9
rect 3 -11 11 9
rect 15 -11 19 9
rect 30 -7 34 13
rect 38 -7 42 13
<< psubstratepcontact >>
rect 30 -47 34 -43
rect -17 -81 -13 -77
rect -8 -81 -4 -77
rect 4 -81 8 -77
rect 15 -81 19 -77
<< nsubstratencontact >>
rect -17 15 -13 19
rect -9 15 -5 19
rect 0 15 4 19
rect 14 15 18 19
rect 30 17 34 22
<< polysilicon >>
rect 35 13 37 16
rect -12 9 -10 12
rect 0 9 2 12
rect 12 9 14 12
rect -12 -41 -10 -11
rect 0 -41 2 -11
rect 12 -41 14 -11
rect 35 -27 37 -7
rect 35 -42 37 -37
rect -12 -75 -10 -71
rect 0 -75 2 -71
rect 12 -75 14 -71
<< polycontact >>
rect -18 -24 -12 -20
rect -6 -31 0 -27
rect 6 -38 12 -34
rect 31 -22 35 -18
<< metal1 >>
rect 30 22 48 23
rect -13 15 -9 19
rect -5 15 0 19
rect 4 15 14 19
rect 18 17 30 19
rect 34 17 48 22
rect 18 15 34 17
rect -17 9 -13 15
rect 3 9 11 15
rect 30 13 34 15
rect -9 -18 -1 -11
rect 15 -18 19 -11
rect 38 -18 42 -7
rect -23 -24 -18 -20
rect -9 -22 31 -18
rect 38 -22 49 -18
rect -23 -31 -6 -27
rect -23 -38 6 -34
rect 15 -41 19 -22
rect 38 -27 42 -22
rect 30 -43 34 -37
rect 34 -47 42 -43
rect -17 -76 -13 -71
rect 30 -76 34 -47
rect -17 -77 34 -76
rect -13 -81 -8 -77
rect -4 -81 4 -77
rect 8 -81 15 -77
rect 19 -81 34 -77
<< labels >>
rlabel metal1 -21 -37 -20 -35 3 a
rlabel metal1 -21 -30 -20 -28 3 b
rlabel metal1 -21 -23 -20 -21 3 c
rlabel metal1 15 -22 19 -18 1 nout
rlabel metal1 -4 -81 4 -76 1 gnd
rlabel ndiffusion -8 -58 -2 -53 1 y
rlabel ndiffusion 4 -58 10 -53 1 x
rlabel metal1 5 14 11 19 1 vdd
rlabel metal1 38 -22 42 -18 1 out
<< end >>
